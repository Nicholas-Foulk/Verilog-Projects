`timescale 1ns / 1ps

module FSM(input [2:0] Op, 
           input Go, clk,
           output [1:0] s1, WA, RAA, RAB, c, s2,
           output WE, REA, REB,
           output [3:0] bcd,
           output DONE
);
  
endmodule
